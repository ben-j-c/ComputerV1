// ClockGenerator.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module ClockGenerator (
		input  wire  ref_clk_clk,        //      ref_clk.clk
		input  wire  ref_reset_reset,    //    ref_reset.reset
		output wire  reset_source_reset, // reset_source.reset
		output wire  sdram_clk_clk,      //    sdram_clk.clk
		output wire  sys_clk_clk         //      sys_clk.clk
	);

	ClockGenerator_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),      //    sdram_clk.clk
		.reset_source_reset (reset_source_reset)  // reset_source.reset
	);

endmodule
