// cordicFixedPoint.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module cordicFixedPoint (
		input  wire [15:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [14:0] c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [14:0] s       //      s.s
	);

	cordicFixedPoint_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
